netcdf \2025-06-16-00.2025-06-17-00.u {
dimensions:
	MT = UNLIMITED ; // (1 currently)
	Y = 3298 ;
	X = 4500 ;
	Depth = 33 ;
variables:
	double MT(MT) ;
		MT:long_name = "time" ;
		MT:units = "days since 1900-12-31 00:00:00" ;
		MT:calendar = "standard" ;
		MT:axis = "T" ;
	double Date(MT) ;
		Date:long_name = "date" ;
		Date:units = "day as %Y%m%d.%f" ;
		Date:C_format = "%13.4f" ;
		Date:FORTRAN_format = "(f13.4)" ;
	float Depth(Depth) ;
		Depth:standard_name = "depth" ;
		Depth:units = "m" ;
		Depth:positive = "down" ;
		Depth:axis = "Z" ;
	int Y(Y) ;
		Y:point_spacing = "even" ;
		Y:axis = "Y" ;
	int X(X) ;
		X:point_spacing = "even" ;
		X:axis = "X" ;
	float Latitude(Y, X) ;
		Latitude:standard_name = "latitude" ;
		Latitude:units = "degrees_north" ;
	float Longitude(Y, X) ;
		Longitude:standard_name = "longitude" ;
		Longitude:units = "degrees_east" ;
		Longitude:modulo = "360 degrees" ;
	float u(MT, Depth, Y, X) ;
		u:coordinates = "Longitude Latitude Date" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:units = "m/s" ;
		u:_FillValue = 1.267651e+30f ;
		u:valid_range = -2.135641f, 2.608399f ;
		u:long_name = " u-veloc. [93.0H]" ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:title = "HYCOM ATLb2.00" ;
		:institution = "National Centers for Environmental Prediction" ;
		:source = "HYCOM archive file" ;
		:experiment = "93.0" ;
		:history = "archv2ncdf3z" ;
}
